/*component round_sig 
	port(
	  ctl : in std_logic;
	  in1 : in std_logic_vector(8 downto 0);
	  values : out std_logic_vector(7 downto 0);
	  back : out std_logic_vector(8 downto 0)
	  );
	end component;

	component round_exp 
	port(
	  ctl : in std_logic;
	  in1 : in std_logic_vector(6 downto 0);
	  values : out std_logic_vector(6 downto 0);
	  back : out std_logic_vector(6 downto 0)
		  );
	end component;*/
